// gps_ca_correlator_channel.sv
// Single-file, Icarus-friendly RTL for one GPS C/A correlator channel with:
//
// Features:
// - Real-only IF input already decoded as fe_val ∈ {+3,+1,-1,-3}
// - GP2021-style 8-phase, 4-level LO (ilo/qlo ∈ {-2,-1,+1,+2})
// - True 0.5-chip Early/Prompt/Late (no dithering)
// - chip_tick aligned to PROMPT chip boundary; dump/epoch counters run on chip_tick
// - Code slew keeps coherent integration length correct by freezing codegen + chip_tick during slewing
// - phase_sync to re-lock half-chip phase convention after slew (safe, non-tick cycle)
//
// NEW in this revision:
// - Adds TIC latch interface (receiver-clock time tag, independent of dump timing)
// - Produces 5 GP2021-like measurement values latched on tic_pulse:
//     TIC_EPOCH
//     TIC_CODE_PHASE (halfchips 0..2046)
//     TIC_CODE_NCO_PHASE (10 MSBs of code NCO accumulator)
//     TIC_CARRIER_CYCLE (20-bit carrier NCO wrap count)
//     TIC_CARRIER_NCO_PHASE (10 MSBs of carrier NCO accumulator)
//
// Notes on code NCO tick:
// - halfchip_tick is generated by MSB edge detect => tick rate is 2 * wrap_rate.
// - If you want nominal halfchip_tick = 2.046 MHz, set code_incr for wrap_rate = 1.023 MHz.
//
// Compile example:
//   iverilog -g2012 -o sim tb.v gps_ca_correlator_channel.sv

`timescale 1ns/1ps

module gps_ca_correlator_channel #(
  parameter integer PHASE_W = 32,
  parameter integer ACC_W   = 18,
  parameter bit     HALFCHIP_OFFSET = 1'b1 // set per your simulator alignment
)(
  input  wire                    clk,
  input  wire                    rstn,

  input  wire                    enable,
  input  wire [7:0]              prn,             // 1..32

  input  wire [31:0]             carr_incr,        // carrier NCO tuning word
  input  wire [31:0]             code_incr,        // code NCO tuning word (see note above)

  input  wire                    slew_req,         // pulse: start slew
  input  wire [10:0]             slew_halfchips,   // number of halfchips to freeze code/dump

  input  wire signed [2:0]       fe_val,           // decoded SIGN/MAG: +/-1 or +/-3

  // TIC: receiver-clock time tag pulse (independent of dump)
  input  wire                    tic_pulse,        // 1clk pulse in SAME clk domain

  output reg                     dump,             // 1clk pulse at end of code period (1023 chips)

  output reg  signed [ACC_W-1:0] i_early,
  output reg  signed [ACC_W-1:0] q_early,
  output reg  signed [ACC_W-1:0] i_prompt,
  output reg  signed [ACC_W-1:0] q_prompt,
  output reg  signed [ACC_W-1:0] i_late,
  output reg  signed [ACC_W-1:0] q_late,

  output reg  [15:0]             code_phase,       // snapshot (chip count 0..1022) at dump
  output reg  [15:0]             carr_phase,       // snapshot (top bits) at dump
  output reg  [15:0]             epoch,            // {unused[15:11], epoch20ms[10:5], epochms[4:0]}
  output reg  [31:0]             dump_count,

  // ---- Measurement registers latched on TIC (GP2021-like) ----
  output reg  [15:0]             tic_epoch,               // epoch sampled at TIC
  output reg  [10:0]             tic_code_phase_halfchip,  // 0..2046 halfchips sampled at TIC
  output reg  [9:0]              tic_code_nco_phase,       // 10 MSBs of code NCO phase accumulator
  output reg  [19:0]             tic_carrier_cycle,        // carrier NCO wrap count sampled at TIC
  output reg  [9:0]              tic_carrier_nco_phase     // 10 MSBs of carrier NCO phase accumulator
);

  // ---------------- Carrier NCO + cycle counter ----------------
  reg  [PHASE_W-1:0] carr_phase_acc;

  // wrap detect using explicit carry-out
  wire [PHASE_W:0] carr_sum  = {1'b0, carr_phase_acc} + {1'b0, carr_incr};
  wire             carr_wrap = carr_sum[PHASE_W]; // 1 when phase wraps: one full 2pi cycle

  always @(posedge clk) begin
    if (!rstn) carr_phase_acc <= {PHASE_W{1'b0}};
    else if (enable) carr_phase_acc <= carr_sum[PHASE_W-1:0];
  end

  // carrier cycle count (20-bit)
  reg [19:0] carrier_cycle_cnt;
  always @(posedge clk) begin
    if (!rstn) carrier_cycle_cnt <= 20'd0;
    else if (enable && carr_wrap) carrier_cycle_cnt <= carrier_cycle_cnt + 20'd1;
  end

  // GP2021-style 8-phase LO, 4-level {-2,-1,+1,+2}
  wire signed [2:0] ilo, qlo;
  carrier_lo_8phase #(.PHASE_W(PHASE_W)) u_lo (
    .phase(carr_phase_acc),
    .ilo(ilo),
    .qlo(qlo)
  );

  // ---------------- Code NCO: half-chip tick via MSB edge ----------------
  reg [PHASE_W-1:0] code_phase_acc;
  reg               code_msb_d;
  wire              halfchip_tick;

  always @(posedge clk) begin
    if (!rstn) begin
      code_phase_acc <= {PHASE_W{1'b0}};
      code_msb_d     <= 1'b0;
    end else if (enable) begin
      code_phase_acc <= code_phase_acc + code_incr;
      code_msb_d     <= code_phase_acc[PHASE_W-1];
    end
  end

  assign halfchip_tick = enable && (code_phase_acc[PHASE_W-1] ^ code_msb_d);

  // ---------------- Slew: freeze codegen and dump timing (coherent length correct) ----------------
  reg        slewing;
  reg [10:0] slew_cnt;

  // countdown in real-time halfchip ticks (fixes off-by-one)
  always @(posedge clk) begin
    if (!rstn) begin
      slewing  <= 1'b0;
      slew_cnt <= 11'd0;
    end else begin
      if (slew_req) begin
        // If 0 requested, do not enter slewing
        slewing  <= (slew_halfchips != 0);
        slew_cnt <= slew_halfchips;
      end

      if (enable && halfchip_tick && slewing) begin
        if (slew_cnt == 11'd1) begin
          // This is the LAST halfchip we want to suppress
          slew_cnt <= 11'd0;
          slewing  <= 1'b0;
        end else begin
          slew_cnt <= slew_cnt - 11'd1;
        end
      end
    end
  end

  // detect slew completion for phase re-lock
  reg slewing_d;
  always @(posedge clk) begin
    if (!rstn) slewing_d <= 1'b0;
    else slewing_d <= slewing;
  end
  wire slew_done = slewing_d && !slewing; // 1-cycle pulse when slewing ends

  // Effective tick that advances code generator (freezes during slew)
  wire halfchip_tick_eff = halfchip_tick && !slewing;

  // ---------------- Code generator: 0.5-chip E/P/L + chip_tick aligned to PROMPT boundary ----------------
  wire ca_e, ca_p, ca_l;
  wire chip_tick;

  // phase_sync: re-lock half_phase to convention after slew (apply only when NOT consuming a tick)
  reg sync_pending;
  always @(posedge clk) begin
    if (!rstn) begin
      sync_pending <= 1'b0;
    end else begin
      if (slew_done) sync_pending <= 1'b1;
      if (phase_sync) sync_pending <= 1'b0;
    end
  end
  wire phase_sync = sync_pending && enable && !halfchip_tick_eff;

  gps_ca_epl_halfchip #(.HALFCHIP_OFFSET(HALFCHIP_OFFSET)) u_ca (
    .clk(clk),
    .rstn(rstn),
    .enable(enable),
    .phase_sync(phase_sync),
    .halfchip_tick(halfchip_tick_eff),
    .prn(prn),
    .early(ca_e),
    .prompt(ca_p),
    .late(ca_l),
    .chip_tick(chip_tick)
  );

  wire signed [1:0] codeE = ca_e ?  2'sd1 : -2'sd1;
  wire signed [1:0] codeP = ca_p ?  2'sd1 : -2'sd1;
  wire signed [1:0] codeL = ca_l ?  2'sd1 : -2'sd1;

  // ---------------- Dump/epoch counters aligned to chip_tick (PROMPT boundary) ----------------
  reg [9:0] chip_cnt; // 0..1022 (1023 chips per code period)

  always @(posedge clk) begin
    if (!rstn) begin
      dump       <= 1'b0;
      dump_count <= 32'd0;
      epoch      <= 16'd0;
      chip_cnt   <= 10'd0;
    end else begin
      dump <= 1'b0;

      if (enable && chip_tick) begin
        if (chip_cnt == 10'd1022) begin
          chip_cnt <= 10'd0;
          dump     <= 1'b1;
          dump_count <= dump_count + 1;

          // epoch[4:0] = 0..19 ms, epoch[10:5] = 0..49 (20ms blocks)
          if (epoch[4:0] == 5'd19) begin
            epoch[4:0] <= 5'd0;
            if (epoch[10:5] == 6'd49) epoch[10:5] <= 6'd0;
            else epoch[10:5] <= epoch[10:5] + 1'b1;
          end else begin
            epoch[4:0] <= epoch[4:0] + 1'b1;
          end
        end else begin
          chip_cnt <= chip_cnt + 1'b1;
        end
      end
    end
  end

  // snapshots for software / logging at dump
  always @(posedge clk) begin
    if (!rstn) begin
      code_phase <= 16'd0;
      carr_phase <= 16'd0;
    end else if (dump) begin
      code_phase <= {6'd0, chip_cnt}; // 0..1022
      carr_phase <= carr_phase_acc[PHASE_W-1 -: 16];
    end
  end

  // ---------------- Continuous CODE_PHASE halfchip counter for TIC ----------------
  // 0..2046, aligned to code generator advancement (frozen during slew)
  reg [10:0] code_halfchip_cnt;
  always @(posedge clk) begin
    if (!rstn) begin
      code_halfchip_cnt <= 11'd0;
    end else if (enable && halfchip_tick_eff) begin
      if (code_halfchip_cnt == 11'd2046)
        code_halfchip_cnt <= 11'd0;
      else
        code_halfchip_cnt <= code_halfchip_cnt + 11'd1;
    end
  end

  // MSBs of NCO accumulators for TIC sampling (GP2021-like)
  wire [9:0] code_nco_phase_msb10_now    = code_phase_acc[PHASE_W-1 -: 10];
  wire [9:0] carrier_nco_phase_msb10_now = carr_phase_acc[PHASE_W-1 -: 10];

  // ---------------- TIC latch: capture 5 measurement values at receiver-clock TIC ----------------
  always @(posedge clk) begin
    if (!rstn) begin
      tic_epoch              <= 16'd0;
      tic_code_phase_halfchip<= 11'd0;
      tic_code_nco_phase     <= 10'd0;
      tic_carrier_cycle      <= 20'd0;
      tic_carrier_nco_phase  <= 10'd0;
    end else if (tic_pulse) begin
      tic_epoch               <= epoch;
      tic_code_phase_halfchip <= code_halfchip_cnt;
      tic_code_nco_phase      <= code_nco_phase_msb10_now;
      tic_carrier_cycle       <= carrier_cycle_cnt;
      tic_carrier_nco_phase   <= carrier_nco_phase_msb10_now;
    end
  end

  // ---------------- Mix ----------------
  // Real input -> complex baseband:
  wire signed [6:0] ibb = fe_val * ilo; // values include 1,2,3,6 (and negative)
  wire signed [6:0] qbb = fe_val * qlo;

  // Code mix for each arm
  wire signed [8:0] ie = ibb * codeE;
  wire signed [8:0] qe = qbb * codeE;
  wire signed [8:0] ip = ibb * codeP;
  wire signed [8:0] qp = qbb * codeP;
  wire signed [8:0] il = ibb * codeL;
  wire signed [8:0] ql = qbb * codeL;

  // ---------------- Accumulate every sample; dump clears ----------------
  reg signed [ACC_W-1:0] acc_ie, acc_qe, acc_ip, acc_qp, acc_il, acc_ql;

  always @(posedge clk) begin
    if (!rstn) begin
      acc_ie <= '0; acc_qe <= '0;
      acc_ip <= '0; acc_qp <= '0;
      acc_il <= '0; acc_ql <= '0;

      i_early  <= '0; q_early  <= '0;
      i_prompt <= '0; q_prompt <= '0;
      i_late   <= '0; q_late   <= '0;
    end else begin
      if (!enable) begin
        acc_ie <= '0; acc_qe <= '0;
        acc_ip <= '0; acc_qp <= '0;
        acc_il <= '0; acc_ql <= '0;
      end else begin
        acc_ie <= acc_ie + {{(ACC_W-9){ie[8]}}, ie};
        acc_qe <= acc_qe + {{(ACC_W-9){qe[8]}}, qe};
        acc_ip <= acc_ip + {{(ACC_W-9){ip[8]}}, ip};
        acc_qp <= acc_qp + {{(ACC_W-9){qp[8]}}, qp};
        acc_il <= acc_il + {{(ACC_W-9){il[8]}}, il};
        acc_ql <= acc_ql + {{(ACC_W-9){ql[8]}}, ql};
      end

      if (dump) begin
        i_early  <= acc_ie; q_early  <= acc_qe;
        i_prompt <= acc_ip; q_prompt <= acc_qp;
        i_late   <= acc_il; q_late   <= acc_ql;

        acc_ie <= '0; acc_qe <= '0;
        acc_ip <= '0; acc_qp <= '0;
        acc_il <= '0; acc_ql <= '0;
      end
    end
  end

endmodule

// ================================================================
// carrier_lo_8phase: GP2021 8-phase, 4-level LO
// ILO: +2 +1 -1 -2 -2 -1 +1 +2 ( cos)
// QLO: -1 -2 -2 -2 +1 +2 +2 +1 (-sin)
// ================================================================
module carrier_lo_8phase #(
  parameter integer PHASE_W = 32
)(
  input  wire [PHASE_W-1:0] phase,
  output reg  signed [2:0]  ilo,
  output reg  signed [2:0]  qlo
);
  wire [2:0] idx = phase[PHASE_W-1 -: 3];

  always @* begin
    case (idx)
      3'd2: begin ilo =  3'sd2; qlo = -3'sd1; end
      3'd3: begin ilo =  3'sd1; qlo = -3'sd2; end
      3'd4: begin ilo = -3'sd1; qlo = -3'sd2; end
      3'd5: begin ilo = -3'sd2; qlo = -3'sd1; end
      3'd6: begin ilo = -3'sd2; qlo =  3'sd1; end
      3'd7: begin ilo = -3'sd1; qlo =  3'sd2; end
      3'd0: begin ilo =  3'sd1; qlo =  3'sd2; end
      3'd1: begin ilo =  3'sd2; qlo =  3'sd1; end
    endcase
  end
endmodule

// ================================================================
// gps_ca_g2_tap_indices: standard GPS L1 C/A PRN 1..32 tap pairs
// ================================================================
module gps_ca_g2_tap_indices(
  input  wire [7:0] prn,
  output reg  [3:0] tapA,
  output reg  [3:0] tapB
);
  always @* begin
    case (prn)
      8'd1:  begin tapA=4'd2; tapB=4'd6;  end
      8'd2:  begin tapA=4'd3; tapB=4'd7;  end
      8'd3:  begin tapA=4'd4; tapB=4'd8;  end
      8'd4:  begin tapA=4'd5; tapB=4'd9;  end
      8'd5:  begin tapA=4'd1; tapB=4'd9;  end
      8'd6:  begin tapA=4'd2; tapB=4'd10; end
      8'd7:  begin tapA=4'd1; tapB=4'd8;  end
      8'd8:  begin tapA=4'd2; tapB=4'd9;  end
      8'd9:  begin tapA=4'd3; tapB=4'd10; end
      8'd10: begin tapA=4'd2; tapB=4'd3;  end
      8'd11: begin tapA=4'd3; tapB=4'd4;  end
      8'd12: begin tapA=4'd5; tapB=4'd6;  end
      8'd13: begin tapA=4'd6; tapB=4'd7;  end
      8'd14: begin tapA=4'd7; tapB=4'd8;  end
      8'd15: begin tapA=4'd8; tapB=4'd9;  end
      8'd16: begin tapA=4'd9; tapB=4'd10; end
      8'd17: begin tapA=4'd1; tapB=4'd4;  end
      8'd18: begin tapA=4'd2; tapB=4'd5;  end
      8'd19: begin tapA=4'd3; tapB=4'd6;  end
      8'd20: begin tapA=4'd4; tapB=4'd7;  end
      8'd21: begin tapA=4'd5; tapB=4'd8;  end
      8'd22: begin tapA=4'd6; tapB=4'd9;  end
      8'd23: begin tapA=4'd1; tapB=4'd3;  end
      8'd24: begin tapA=4'd4; tapB=4'd6;  end
      8'd25: begin tapA=4'd5; tapB=4'd7;  end
      8'd26: begin tapA=4'd6; tapB=4'd8;  end
      8'd27: begin tapA=4'd7; tapB=4'd9;  end
      8'd28: begin tapA=4'd8; tapB=4'd10; end
      8'd29: begin tapA=4'd1; tapB=4'd6;  end
      8'd30: begin tapA=4'd2; tapB=4'd7;  end
      8'd31: begin tapA=4'd3; tapB=4'd8;  end
      8'd32: begin tapA=4'd4; tapB=4'd9;  end
      default: begin tapA=4'd2; tapB=4'd6; end
    endcase
  end
endmodule

// ================================================================
// gps_ca_epl_halfchip: true 0.5-chip Early/Prompt/Late
// - phase_sync re-locks half_phase to HALFCHIP_OFFSET without resetting LFSRs,
//   preventing half-chip convention flips after slew.
// - chip_tick pulses on second half of each chip (aligned to PROMPT chip boundary).
// ================================================================
module gps_ca_epl_halfchip #(
  parameter bit HALFCHIP_OFFSET = 1'b0
)(
  input  wire       clk,
  input  wire       rstn,
  input  wire       enable,
  input  wire       phase_sync,
  input  wire       halfchip_tick,
  input  wire [7:0] prn,

  output reg        early,
  output reg        prompt,
  output reg        late,
  output wire       chip_tick
);
  reg [9:0] g1, g2;
  reg       half_phase; // 0 first half, 1 second half

  wire [3:0] tapA, tapB;
  gps_ca_g2_tap_indices u_idx(.prn(prn), .tapA(tapA), .tapB(tapB));

  function automatic bit pick_stage(input [9:0] s, input [3:0] pos1b);
    begin
      pick_stage = s[pos1b-1];
    end
  endfunction

  // current chip from current states
  wire g1_out = g1[9];
  wire g2_out = pick_stage(g2, tapA) ^ pick_stage(g2, tapB);
  wire chip_curr = g1_out ^ g2_out;

  // feedback polynomials
  wire g1_fb = g1[2] ^ g1[9];
  wire g2_fb = g2[1] ^ g2[2] ^ g2[5] ^ g2[7] ^ g2[8] ^ g2[9];

  // next states / next chip for +0.5-chip late on second half
  wire [9:0] g1_next = {g1[8:0], g1_fb};
  wire [9:0] g2_next = {g2[8:0], g2_fb};
  wire chip_next = g1_next[9] ^ (pick_stage(g2_next, tapA) ^ pick_stage(g2_next, tapB));

  reg chip_prev;

  // Chip tick aligned to PROMPT boundary: pulse on second half of each chip
  assign chip_tick = enable && halfchip_tick && (half_phase == 1'b1);

  always @(posedge clk) begin
    if (!rstn) begin
      g1 <= 10'h3FF;
      g2 <= 10'h3FF;
      half_phase <= HALFCHIP_OFFSET;
      chip_prev  <= 1'b1;
      early <= 1'b1; prompt <= 1'b1; late <= 1'b1;
    end else begin
      if (phase_sync) begin
        // Re-lock half-chip convention safely on a non-tick cycle
        half_phase <= HALFCHIP_OFFSET;
      end else if (enable && halfchip_tick) begin
        // 0.5-chip E/P/L:
        if (!half_phase) begin
          early  <= chip_prev;
          prompt <= chip_curr;
          late   <= chip_curr;
        end else begin
          early  <= chip_curr;
          prompt <= chip_curr;
          late   <= chip_next;
        end

        // advance LFSRs on chip boundary (after second half)
        if (half_phase) begin
          g1 <= g1_next;
          g2 <= g2_next;
          chip_prev <= chip_curr;
        end

        half_phase <= ~half_phase;
      end
    end
  end
endmodule
